//------------------------------------------------------------------------------------------------------------------//
// FILE NAME       : apb_i2c_defines.sv 
// AUTHOR          : Harekrishna ray
// MODIFIED DATE   : 20/02/23
// DESCRIPTION     : file contains the different defines 
//------------------------------------------------------------------------------------------------------------------//


`define ADDR_WIDTH 8
`define DATA_WIDTH 8

`define DEPTH 8
